module song_rom (	input clk,				
	input [6:0] addr,				
	output reg [15:0] dout				
					
);					
	wire [15:0] memory [127:0];				
					
	always @(posedge clk)				
		dout = memory[addr];			
					
	assign memory[	  0	] =	{1'b0, 6'd40, 6'd48, 3'd0};	// Note: 4C
	assign memory[	  1	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	  2	] =	{1'b0, 6'd44, 6'd36, 3'd0};	// Note: 4E
	assign memory[	  3	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	  4	] =	{1'b0, 6'd47, 6'd24, 3'd0};	// Note: 4G
	assign memory[	  5	] =	{1'd1, 6'd24, 9'd0};	// Note: 
	assign memory[	  6	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	  7	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	  8	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	  9	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 10	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 11	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 12	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 13	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 14	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 15	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 16	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 17	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 18	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 19	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 20	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 21	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 22	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 23	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 24	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 25	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 26	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 27	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 28	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 29	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 30	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 31	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 32	] =	{1'b0, 6'd40, 6'd12, 3'd0};	// Note: 4C
	assign memory[	 33	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 34	] =	{1'b0, 6'd41, 6'd12, 3'd0};	// Note: 4C#Db
	assign memory[	 35	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 36	] =	{1'b0, 6'd42, 6'd12, 3'd0};	// Note: 4D
	assign memory[	 37	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 38	] =	{1'b0, 6'd43, 6'd12, 3'd0};	// Note: 4D#Eb
	assign memory[	 39	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 40	] =	{1'b0, 6'd44, 6'd12, 3'd0};	// Note: 4E
	assign memory[	 41	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 42	] =	{1'b0, 6'd45, 6'd12, 3'd0};	// Note: 4F
	assign memory[	 43	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 44	] =	{1'b0, 6'd46, 6'd12, 3'd0};	// Note: 4F#Gb
	assign memory[	 45	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 46	] =	{1'b0, 6'd47, 6'd12, 3'd0};	// Note: 4G
	assign memory[	 47	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 48	] =	{1'b0, 6'd48, 6'd12, 3'd0};	// Note: 4G#Ab
	assign memory[	 49	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 50	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 51	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 52	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 53	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 54	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 55	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 56	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 57	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 58	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 59	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 60	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 61	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 62	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 63	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 64	] =	{1'b0, 6'd52, 6'd48, 3'd0};	// Note: 5C
	assign memory[	 65	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 66	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 67	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 68	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 69	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 70	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 71	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 72	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 73	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 74	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 75	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 76	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 77	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 78	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 79	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 80	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 81	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 82	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 83	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 84	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 85	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 86	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 87	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 88	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 89	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 90	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 91	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 92	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 93	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 94	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 95	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 96	] =	{1'b0, 6'd40, 6'd48, 3'd0};	// Note: 4C
	assign memory[	 97	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 98	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 99	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	100	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	101	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	102	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	103	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	104	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	105	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	106	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	107	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	108	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	109	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	110	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	111	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	112	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	113	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	114	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	115	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	116	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	117	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	118	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	119	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	120	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	121	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	122	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	123	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	124	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	125	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	126	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	127	] =	{1'd1, 6'd0, 9'd0};	// Note: 
					
endmodule					
