module song_rom5 (	input clk,				
	input [8:0] addr,				
	output reg [15:0] dout				
					
);					
	wire [15:0] memory [511:0];				
					
	always @(posedge clk)				
		dout = memory[addr];			
					
	assign memory[	  0	] =	{1'b0, 6'd11, 6'd12, 3'd0};	// Note: 1G
	assign memory[	  1	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	  2	] =	{1'b0, 6'd11, 6'd12, 3'd0};	// Note: 1G
	assign memory[	  3	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	  4	] =	{1'b0, 6'd11, 6'd12, 3'd0};	// Note: 1G
	assign memory[	  5	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	  6	] =	{1'b0, 6'd11, 6'd12, 3'd0};	// Note: 1G
	assign memory[	  7	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	  8	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	  9	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 10	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 11	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 12	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 13	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 14	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 15	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 16	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 17	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 18	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 19	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 20	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 21	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 22	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 23	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 24	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 25	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 26	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 27	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 28	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 29	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 30	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 31	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 32	] =	{1'b0, 6'd11, 6'd12, 3'd0};	// Note: 1G
	assign memory[	 33	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 34	] =	{1'b0, 6'd14, 6'd12, 3'd0};	// Note: 2A#Bb
	assign memory[	 35	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 36	] =	{1'b0, 6'd16, 6'd12, 3'd0};	// Note: 2C
	assign memory[	 37	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 38	] =	{1'b0, 6'd14, 6'd12, 3'd0};	// Note: 2A#Bb
	assign memory[	 39	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 40	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	 41	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 42	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	 43	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 44	] =	{1'b0, 6'd28, 6'd12, 3'd0};	// Note: 3C
	assign memory[	 45	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 46	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	 47	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 48	] =	{1'b0, 6'd30, 6'd12, 3'd0};	// Note: 3D
	assign memory[	 49	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 50	] =	{1'b0, 6'd28, 6'd12, 3'd0};	// Note: 3C
	assign memory[	 51	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 52	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	 53	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 54	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	 55	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 56	] =	{1'b0, 6'd21, 6'd12, 3'd0};	// Note: 2F
	assign memory[	 57	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 58	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	 59	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 60	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	 61	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 62	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	 63	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 64	] =	{1'b0, 6'd38, 6'd12, 3'd0};	// Note: 4A#Bb
	assign memory[	 65	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 66	] =	{1'b0, 6'd38, 6'd12, 3'd0};	// Note: 4A#Bb
	assign memory[	 67	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 68	] =	{1'b0, 6'd35, 6'd12, 3'd0};	// Note: 3G
	assign memory[	 69	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 70	] =	{1'b0, 6'd35, 6'd12, 3'd0};	// Note: 3G
	assign memory[	 71	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 72	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 73	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 74	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 75	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 76	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 77	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 78	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 79	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 80	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 81	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 82	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 83	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 84	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 85	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 86	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 87	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 88	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 89	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 90	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 91	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 92	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 93	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 94	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 95	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	 96	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	 97	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	 98	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	 99	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	100	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	101	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	102	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	103	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	104	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	105	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	106	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	107	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	108	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	109	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	110	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	111	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	112	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	113	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	114	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	115	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	116	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	117	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	118	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	119	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	120	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	121	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	122	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	123	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	124	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	125	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	126	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	127	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	128	] =	{1'b0, 6'd21, 6'd12, 3'd0};	// Note: 2F
	assign memory[	129	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	130	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	131	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	132	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	133	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	134	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	135	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	136	] =	{1'b0, 6'd30, 6'd12, 3'd0};	// Note: 3D
	assign memory[	137	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	138	] =	{1'b0, 6'd23, 6'd6, 3'd0};	// Note: 2G
	assign memory[	139	] =	{1'd1, 6'd6, 9'd0};	// Note: 
	assign memory[	140	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	141	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	142	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	143	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	144	] =	{1'b0, 6'd21, 6'd18, 3'd0};	// Note: 2F
	assign memory[	145	] =	{1'd1, 6'd18, 9'd0};	// Note: 
	assign memory[	146	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	147	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	148	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	149	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	150	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	151	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	152	] =	{1'b0, 6'd30, 6'd12, 3'd0};	// Note: 3D
	assign memory[	153	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	154	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	155	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	156	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	157	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	158	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	159	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	160	] =	{1'b0, 6'd11, 6'd12, 3'd0};	// Note: 1G
	assign memory[	161	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	162	] =	{1'b0, 6'd14, 6'd12, 3'd0};	// Note: 2A#Bb
	assign memory[	163	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	164	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	165	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	166	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	167	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	168	] =	{1'b0, 6'd30, 6'd12, 3'd0};	// Note: 3D
	assign memory[	169	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	170	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	171	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	172	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	173	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	174	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	175	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	176	] =	{1'b0, 6'd9, 6'd12, 3'd0};	// Note: 1F
	assign memory[	177	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	178	] =	{1'b0, 6'd21, 6'd12, 3'd0};	// Note: 2F
	assign memory[	179	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	180	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	181	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	182	] =	{1'b0, 6'd21, 6'd12, 3'd0};	// Note: 2F
	assign memory[	183	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	184	] =	{1'b0, 6'd28, 6'd12, 3'd0};	// Note: 3C
	assign memory[	185	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	186	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	187	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	188	] =	{1'b0, 6'd25, 6'd12, 3'd0};	// Note: 3A
	assign memory[	189	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	190	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	191	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	192	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	193	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	194	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	195	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	196	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	197	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	198	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	199	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	200	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	201	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	202	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	203	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	204	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	205	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	206	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	207	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	208	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	209	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	210	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	211	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	212	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	213	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	214	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	215	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	216	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	217	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	218	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	219	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	220	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	221	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	222	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	223	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	224	] =	{1'b0, 6'd21, 6'd6, 3'd0};	// Note: 2F
	assign memory[	225	] =	{1'd1, 6'd6, 9'd0};	// Note: 
	assign memory[	226	] =	{1'b0, 6'd23, 6'd6, 3'd0};	// Note: 2G
	assign memory[	227	] =	{1'd1, 6'd6, 9'd0};	// Note: 
	assign memory[	228	] =	{1'b0, 6'd26, 6'd6, 3'd0};	// Note: 3A#Bb
	assign memory[	229	] =	{1'd1, 6'd6, 9'd0};	// Note: 
	assign memory[	230	] =	{1'b0, 6'd28, 6'd12, 3'd0};	// Note: 3C
	assign memory[	231	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	232	] =	{1'b0, 6'd26, 6'd6, 3'd0};	// Note: 3A#Bb
	assign memory[	233	] =	{1'd1, 6'd6, 9'd0};	// Note: 
	assign memory[	234	] =	{1'b0, 6'd30, 6'd12, 3'd0};	// Note: 3D
	assign memory[	235	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	236	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	237	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	238	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	239	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	240	] =	{1'b0, 6'd21, 6'd12, 3'd0};	// Note: 2F
	assign memory[	241	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	242	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	243	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	244	] =	{1'b0, 6'd16, 6'd12, 3'd0};	// Note: 2C
	assign memory[	245	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	246	] =	{1'b0, 6'd18, 6'd12, 3'd0};	// Note: 2D
	assign memory[	247	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	248	] =	{1'b0, 6'd23, 6'd12, 3'd0};	// Note: 2G
	assign memory[	249	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	250	] =	{1'b0, 6'd26, 6'd12, 3'd0};	// Note: 3A#Bb
	assign memory[	251	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	252	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	253	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	254	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	255	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	256	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	257	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	258	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	259	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	260	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	261	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	262	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	263	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	264	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	265	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	266	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	267	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	268	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	269	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	270	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	271	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	272	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	273	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	274	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	275	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	276	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	277	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	278	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	279	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	280	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	281	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	282	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	283	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	284	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	285	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	286	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	287	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	288	] =	{1'b0, 6'd19, 6'd12, 3'd0};	// Note: 2D#Eb
	assign memory[	289	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	290	] =	{1'b0, 6'd31, 6'd12, 3'd0};	// Note: 3D#Eb
	assign memory[	291	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	292	] =	{1'b0, 6'd35, 6'd12, 3'd0};	// Note: 3G
	assign memory[	293	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	294	] =	{1'b0, 6'd31, 6'd12, 3'd0};	// Note: 3D#Eb
	assign memory[	295	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	296	] =	{1'b0, 6'd40, 6'd12, 3'd0};	// Note: 4C
	assign memory[	297	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	298	] =	{1'b0, 6'd38, 6'd12, 3'd0};	// Note: 4A#Bb
	assign memory[	299	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	300	] =	{1'b0, 6'd35, 6'd12, 3'd0};	// Note: 3G
	assign memory[	301	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	302	] =	{1'b0, 6'd31, 6'd12, 3'd0};	// Note: 3D#Eb
	assign memory[	303	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	304	] =	{1'b0, 6'd31, 6'd12, 3'd0};	// Note: 3D#Eb
	assign memory[	305	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	306	] =	{1'b0, 6'd31, 6'd12, 3'd0};	// Note: 3D#Eb
	assign memory[	307	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	308	] =	{1'b0, 6'd35, 6'd12, 3'd0};	// Note: 3G
	assign memory[	309	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	310	] =	{1'b0, 6'd38, 6'd12, 3'd0};	// Note: 4A#Bb
	assign memory[	311	] =	{1'd1, 6'd12, 9'd0};	// Note: 
	assign memory[	312	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	313	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	314	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	315	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	316	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	317	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	318	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	319	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	320	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	321	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	322	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	323	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	324	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	325	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	326	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	327	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	328	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	329	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	330	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	331	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	332	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	333	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	334	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	335	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	336	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	337	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	338	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	339	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	340	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	341	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	342	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	343	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	344	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	345	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	346	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	347	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	348	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	349	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	350	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	351	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	352	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	353	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	354	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	355	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	356	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	357	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	358	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	359	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	360	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	361	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	362	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	363	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	364	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	365	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	366	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	367	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	368	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	369	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	370	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	371	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	372	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	373	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	374	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	375	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	376	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	377	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	378	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	379	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	380	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	381	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	382	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	383	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	384	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	385	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	386	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	387	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	388	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	389	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	390	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	391	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	392	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	393	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	394	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	395	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	396	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	397	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	398	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	399	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	400	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	401	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	402	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	403	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	404	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	405	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	406	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	407	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	408	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	409	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	410	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	411	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	412	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	413	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	414	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	415	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	416	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	417	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	418	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	419	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	420	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	421	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	422	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	423	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	424	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	425	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	426	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	427	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	428	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	429	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	430	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	431	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	432	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	433	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	434	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	435	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	436	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	437	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	438	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	439	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	440	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	441	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	442	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	443	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	444	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	445	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	446	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	447	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	448	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	449	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	450	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	451	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	452	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	453	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	454	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	455	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	456	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	457	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	458	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	459	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	460	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	461	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	462	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	463	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	464	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	465	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	466	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	467	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	468	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	469	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	470	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	471	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	472	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	473	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	474	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	475	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	476	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	477	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	478	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	479	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	480	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	481	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	482	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	483	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	484	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	485	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	486	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	487	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	488	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	489	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	490	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	491	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	492	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	493	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	494	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	495	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	496	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	497	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	498	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	499	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	500	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	501	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	502	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	503	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	504	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	505	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	506	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	507	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	508	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	509	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	510	] =	{1'd1, 6'd0, 9'd0};	// Note: 
	assign memory[	511	] =	{1'd1, 6'd0, 9'd0};	// Note: 
					
endmodule					