/* SKELETON CODE
* module distributor */
